module compute_tb ();

endmodule
