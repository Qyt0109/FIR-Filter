module delay_pipeline_tb ();

endmodule
