module filter_tb ();

endmodule
