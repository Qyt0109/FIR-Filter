module coeffs ();

endmodule
