module counter #(
    parameter MAX_COUNT = 100
) (
    input clk
);

endmodule
