module counter_tb ();

endmodule
