module delay_pipeline ();

endmodule
