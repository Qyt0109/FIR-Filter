module filter ();

endmodule
