module compute ();

endmodule
